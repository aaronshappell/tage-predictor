`ifndef COMMON_DEFINES_SVH
`define COMMON_DEFINES_SVH

`define BR_TAKEN        1'b1
`define BR_NOT_TAKEN    1'b0

`define BHT_IDX_WIDTH   11
`define TAGE_IDX_WIDTH  `BHT_IDX_WIDTH - 2

`endif