`include "common_defines.svh"

module tage_predictor
    (
        input logic clk_i,
        input logic [`TAGE_IDX_WIDTH-1:0] w_idx_i,
        input logic br_result_i,
        input logic [`TAGE_IDX_WIDTH-1:0] r_idx_i,
        output logic prediction_o
    );

endmodule
