`ifndef COMMON_DEFINES_SVH
`define COMMON_DEFINES_SVH

`define BR_TAKEN        1'b1
`define BR_NOT_TAKEN    1'b0

`define IDX_WIDTH       9

`endif